library verilog;
use verilog.vl_types.all;
entity my_dff_vlg_sample_tst is
    port(
        C               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end my_dff_vlg_sample_tst;
