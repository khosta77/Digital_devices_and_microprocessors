library verilog;
use verilog.vl_types.all;
entity decoder_20L274_vlg_vec_tst is
end decoder_20L274_vlg_vec_tst;
