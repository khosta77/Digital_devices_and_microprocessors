library verilog;
use verilog.vl_types.all;
entity two_circuit_vlg_vec_tst is
end two_circuit_vlg_vec_tst;
