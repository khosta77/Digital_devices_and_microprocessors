library verilog;
use verilog.vl_types.all;
entity VD2_20_vlg_vec_tst is
end VD2_20_vlg_vec_tst;
