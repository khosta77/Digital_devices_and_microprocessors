library verilog;
use verilog.vl_types.all;
entity bsd_vlg_vec_tst is
end bsd_vlg_vec_tst;
