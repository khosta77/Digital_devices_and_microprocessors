library verilog;
use verilog.vl_types.all;
entity VD2_20_vlg_sample_tst is
    port(
        START           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end VD2_20_vlg_sample_tst;
