library verilog;
use verilog.vl_types.all;
entity VD2_20 is
    port(
        \OUT\           : out    vl_logic;
        \IN\            : in     vl_logic
    );
end VD2_20;
