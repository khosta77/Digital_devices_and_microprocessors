library verilog;
use verilog.vl_types.all;
entity CNT_vlg_vec_tst is
end CNT_vlg_vec_tst;
