library verilog;
use verilog.vl_types.all;
entity asynchronous_counter_vlg_vec_tst is
end asynchronous_counter_vlg_vec_tst;
