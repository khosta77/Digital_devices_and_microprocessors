library verilog;
use verilog.vl_types.all;
entity \2_circuit\ is
    port(
        A1              : out    vl_logic;
        X3              : in     vl_logic;
        X2              : in     vl_logic;
        X1              : in     vl_logic;
        X0              : in     vl_logic
    );
end \2_circuit\;
