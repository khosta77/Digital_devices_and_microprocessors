library verilog;
use verilog.vl_types.all;
entity VD2_20_vlg_check_tst is
    port(
        \OUT\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end VD2_20_vlg_check_tst;
