library verilog;
use verilog.vl_types.all;
entity decoder_20L274 is
    port(
        X0              : out    vl_logic;
        A2              : in     vl_logic;
        A1              : in     vl_logic;
        A0              : in     vl_logic;
        X1              : out    vl_logic;
        X2              : out    vl_logic;
        X3              : out    vl_logic
    );
end decoder_20L274;
