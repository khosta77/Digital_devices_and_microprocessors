library verilog;
use verilog.vl_types.all;
entity decoder_20L274_vlg_check_tst is
    port(
        X0              : in     vl_logic;
        X1              : in     vl_logic;
        X2              : in     vl_logic;
        X3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder_20L274_vlg_check_tst;
