library verilog;
use verilog.vl_types.all;
entity my_dff_vlg_vec_tst is
end my_dff_vlg_vec_tst;
